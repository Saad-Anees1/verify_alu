class alu_seqr extends uvm_sequencer #(alu_seq_item);
  `uvm_component_utils(alu_seqr)

 `uvm_component_new

endclass
