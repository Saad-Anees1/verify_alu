package alu_pkg;
  import uvm_pkg::*;
  import alu_types_pkg::*;

  `include "uvm_macros.svh"
  `include "dv_macros.svh"

  `include "alu_seq_item.sv"
  `include "alu_env_cfg.sv"
  `include "alu_seq.sv"
  `include "div0_seq_c.sv"
  `include "alu_add.sv"
  `include "alu_sub.sv"
  `include "alu_nop.sv"
  `include "alu_seqr.sv"
  `include "alu_drv.sv"
  `include "alu_mon.sv"
  `include "alu_agent.sv"
  `include "alu_scb.sv"
  `include "alu_coverage.sv"
  `include "alu_env.sv"
  `include "alu_test.sv"

endpackage
