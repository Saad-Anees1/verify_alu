class div0_seq_c extends alu_seq;
  `uvm_object_utils(div0_seq_c)

  `uvm_object_new

  task body();
    $display("calling div0_seq_c seq....");
  endtask
endclass
